    bbb1100qweex0 wertx0 ertex00rtyex0(x=3;x++;x++;x--;!a5;!b3;!c5;end;x=3;x++;x++;x--;!a5;!b3;!c5;end;x=3;x++;!a3;!a3;!b3;!c2;x++;x++;x++;x++;x++;end;x=3;x++;x++;x++;!a2;!a1;!b2;!c1;!a2;end;