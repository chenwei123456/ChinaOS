     aaa1100aaa1100cccex0i=9;i++;end;